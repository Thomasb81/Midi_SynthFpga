`timescale 1ns / 1ps
module event_48k_gene(
    input clk,
    input rst,
    output [47:0] events
    );

reg [9:0] count;

always @(posedge clk)
if (rst==1'b1)
  count <= 10'h000;
else if (count == 666)
  count <= 10'h000;
else
  count <= count + 1;

assign events = 
(count == 0  ) ? 48'h000000000001 :
(count == 1  ) ? 48'h000000000002 :
(count == 2  ) ? 48'h000000000004 :
(count == 3  ) ? 48'h000000000008 :
(count == 4  ) ? 48'h000000000010 :
(count == 5  ) ? 48'h000000000020 :
(count == 6  ) ? 48'h000000000040 :
(count == 7  ) ? 48'h000000000080 :
(count == 8  ) ? 48'h000000000100 :
(count == 9  ) ? 48'h000000000200 :
(count == 10 ) ? 48'h000000000400 :
(count == 11 ) ? 48'h000000000800 :
(count == 12 ) ? 48'h000000001000 :
(count == 13 ) ? 48'h000000002000 :
(count == 14 ) ? 48'h000000004000 :
(count == 15 ) ? 48'h000000008000 :
(count == 16 ) ? 48'h000000010000 :
(count == 17 ) ? 48'h000000020000 :
(count == 18 ) ? 48'h000000040000 :
(count == 19 ) ? 48'h000000080000 :
(count == 20 ) ? 48'h000000100000 :
(count == 21 ) ? 48'h000000200000 :
(count == 22 ) ? 48'h000000400000 :
(count == 23 ) ? 48'h000000800000 :
(count == 24 ) ? 48'h000001000000 :
(count == 25 ) ? 48'h000002000000 :
(count == 26 ) ? 48'h000004000000 :
(count == 27 ) ? 48'h000008000000 :
(count == 28 ) ? 48'h000010000000 :
(count == 29 ) ? 48'h000020000000 :
(count == 30 ) ? 48'h000040000000 :
(count == 31 ) ? 48'h000080000000 :
(count == 32 ) ? 48'h000100000000 :
(count == 33 ) ? 48'h000200000000 :
(count == 34 ) ? 48'h000400000000 :
(count == 35 ) ? 48'h000800000000 :
(count == 36 ) ? 48'h001000000000 :
(count == 37 ) ? 48'h002000000000 :
(count == 38 ) ? 48'h004000000000 :
(count == 39 ) ? 48'h008000000000 :
(count == 40 ) ? 48'h010000000000 :
(count == 41 ) ? 48'h020000000000 :
(count == 42 ) ? 48'h040000000000 :
(count == 43 ) ? 48'h080000000000 :
(count == 44 ) ? 48'h100000000000 :
(count == 45 ) ? 48'h200000000000 :
(count == 46 ) ? 48'h400000000000 :
(count == 47 ) ? 48'h800000000000 :
48'h0000000000;

endmodule
