
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library UNISIM;
use UNISIM.VComponents.all;


entity RAMB16_S18_wavetable is
  Port (clk : in std_logic;
        addr : in std_logic_vector (9 downto 0);
        en : in std_logic;
        do : out std_logic_vector (17 downto 0)
       );
end RAMB16_S18_wavetable;

architecture Behav of RAMB16_S18_wavetable is


begin

RAMB16_S18_inst0 : RAMB16_S18
   generic map (
      INIT => X"000",
      SRVAL => X"000",
      INIT_00 => X"689d69d76acb6b596b706b0b6a336901679d663464fa641e63cc6422652c66e6",
      INIT_01 => X"7b12786a759372a36fb36ce06a4567fe662564ce640363c9641764da65f56744",
      INIT_02 => X"7699785c7a3c7c267e057fc18145827e835c83d183d8836c828e81417f8c7d78",
      INIT_03 => X"623063c36574672e68da6a686bcb6cfe6e056ee86fb970887169726c739c7501",
      INIT_04 => X"4bd94f13522854f65762595d5ae15bf65cae5d235d765dc75e325ed05fad60cf",
      INIT_05 => X"1fe323ea27d82b822eca31a43414362c380c39d63baf3db74002429b457f489c",
      INIT_06 => X"156917cb191b196518cb178415d81416128c1180112c11b0131b156218661bf9",
      INIT_07 => X"da58ddffe0e9e350e577e7a2ea13ecfbf079f498f948fe6303b008ea0dc91206",
      INIT_08 => X"70fd746278657d2182a98905902c9804a064a914b1d3ba5dc26dc9cad047d5cc",
      INIT_09 => X"4df5506352a554c756d458d75ad75cd95ede60e662f064fd6712693b6b896e15",
      INIT_0A => X"1f3b20a822702490270329c72cd5302233a0373c3ae33e804201455448714b51",
      INIT_0B => X"652e5b18515148103f8437d731232b7926dc2343209c1ed21dc71d631d8c1e2e",
      INIT_0C => X"d4adcffdcb46c681c19fbc8cb732b178ab44a4819d1d95128c63832179666f5a",
      INIT_0D => X"224a1d64185c13450e2d091e0421ff37fa5ff597f0daec24e771e2bfde0dd95d",
      INIT_0E => X"4f8a4d7b4b654952474745414337411c3edf3c6e39b936b0334d2f8a2b6d26fd",
      INIT_0F => X"512f52c0541c554b5653573157e2585d589758875824576b565c54fe535d5186",
      INIT_10 => X"1d0d1f4821f5251228992c78309634d439133d33411a44b247ed4ac64d3e4f5d",
      INIT_11 => X"13c112a511dc1171116211a7123012e813be14a2158a1677176e187e19ba1b38",
      INIT_12 => X"11ed119b1206130b147b161e17be19261a2d1ab81abb1a3b194918041692151a",
      INIT_13 => X"2d582e302ef22f6d2f732edd2d942b9228e525ad221b1e6a1ad717a014fb130d",
      INIT_14 => X"1fe323d327622a602cb02e402f162f442eef2e452d782cb82c2f2bf82c1e2c9c",
      INIT_15 => X"03050443054d061a06ae0719077907f308ad09ce0b740db1108713e817b71bc7",
      INIT_16 => X"fe12ff7d005e00b4008d0005ff43fe71fdb9fd3ffd1efd62fe0cff0c004a01a8",
      INIT_17 => X"f009f0dcf10af0bbf021ef74eeebeeb5eef6efc2f11bf2f1f524f78af9f3fc2f",
      INIT_18 => X"af27b3c4b829bc6dc0a9c4f5c965ce00d2c2d799dc66e105e548e907ec1fee78",
      INIT_19 => X"8fcc8c3988f38646847383a98405858c88308bcd903295279a6f9fd4a527aa48",
      INIT_1A => X"7dd9814084eb88c28ca690739401972499ae9b779c5e9c4f9b49995996a5935f",
      INIT_1B => X"bb52afdba4b69a4090cb889181ba7c55785e75c27461741574b7762178327acd",
      INIT_1C => X"08b8056202d500feffb1feadfd9dfc27f9eff6a5f20dec02e480dba0d197c6b3",
      INIT_1D => X"438e3fd33cc53a41381135f933ba311c2df72a3725dd21041bd81695117c0ccb",
      INIT_1E => X"6faa71cc73c17544761175ef74b672536ecf6a4764ef5f0e58ef52e14d2b4804",
      INIT_1F => X"69976a866b606c066c606c646c166b876ad56a2769a5697869bf6a8a6bda6d9c",
      INIT_20 => X"718d71ef71f8719d70df6fc86e6e6ced6b6769ff68d76806679d679e680368b4",
      INIT_21 => X"7924773f7553737571b7702c6ee46dee6d526d146d326da16e506f28700e70e4",
      INIT_22 => X"761877b379517ae77c677dc17ee77fc9805b809680757ff97f247dff7c947af1",
      INIT_23 => X"51d053f8568d59705c7d5f91628e655d67ee6a3c6c4a6e226fd2716972f67483",
      INIT_24 => X"3b463faf43e447a94ace4d364ed64fb94ffb4fc84f544ed84e894e944f1a502d",
      INIT_25 => X"25292792295e2a7b2aef2ad52a5b29bb2937290f297c2aa52c9e2f6532e336ec",
      INIT_26 => X"12d9149e157f159d152b146a139e130c12ee136e14a2168819091bfa1f242249",
      INIT_27 => X"d572d85adaf3dd71e009e2ede642ea1fee86f367f89ffdfd034208310c8d1025",
      INIT_28 => X"78e67d4e823487a08d8f93f99acaa1e4a920b053b74ebde5c3f1c958ce0bd20e",
      INIT_29 => X"4b6e4e41510153ad564858d55b585dd8605a62e5658068336b0a6e11715874ee",
      INIT_2A => X"238b25d028092a332c512e6c309032c8351c37943a2f3cec3fc442ac459d488a",
      INIT_2B => X"58534df043fe3ac032702b41255520bd1d7b1b7c1aa31ac51bb21d361f212149",
      INIT_2C => X"d285cce2c731c175bba6b5b9af97a929a2549afe93128a85815777976d6262e4",
      INIT_2D => X"1af3169912540e280a160616021efe1ffa0cf5d3f16aecc8e7ebe2d3dd89d816",
      INIT_2E => X"4902480f46e7458643e642013fd23d553a85376333f130352c3a280c23bb1f59",
      INIT_2F => X"4f424ee04e5d4dcf4d444cca4c654c174bde4bb14b8a4b5e4b234ad04a5e49c6",
      INIT_30 => X"298b2ca63006339b374f3b0b3eb4422d455f48314a944c7b4de44ed34f514f70",
      INIT_31 => X"1efe1ed31e7a1e091d951d301cec1cd71cfd1d661e1c1f232081223a244f26c1",
      INIT_32 => X"159f138612071134110f118e129b141615d717b819911b411cae1dc71e851ee9",
      INIT_33 => X"2b942ada2a802a6f2a882aa32a932a322960280b262d23d421171e1f1b171832",
      INIT_34 => X"139819441f00247f29782db130fc3342348034c8343e331631872fcf2e232cb0",
      INIT_35 => X"065f06a8068905fe051003d7027b012b0020ff93ffb900ba02b105a7098e0e45",
      INIT_36 => X"003a0105017d01aa019c0167012500f100e2010a0172021802f203e904e305bf",
      INIT_37 => X"f03ff0e3f151f1a1f1ecf249f2cdf388f482f5bdf730f8cdfa7ffc2dfdc0ff20",
      INIT_38 => X"b794bcd9c21ac744cc47d116d5a8d9f3ddf1e19ae4e5e7cdea4dec61ee0cef52",
      INIT_39 => X"a686a425a19f9f2a9cfb9b439a2c99d69a539bad9ddda0d5a47ea8b9ad66b265",
      INIT_3A => X"865c89e38da89197959b99999d76a112a44ba702a91aaa7cab1caaf6aa15a88f",
      INIT_3B => X"b440aa43a0c6980c904d89b1844f802f7d4a7b8f7ae37b277c3a7dfe80558326",
      INIT_3C => X"0fc00c390913063a038700c8fdc3fa3bf5f9f0d2eaa9e377db47d23cc88abe72",
      INIT_3D => X"42a93fb33d503b57399437d135db338830bd2d6e29a3257020fa1c6b17ee13ac",
      INIT_3E => X"6e197104735174c37529746372696f466b1d6624609d5ad455114f984aa0464b",
      INIT_3F => X"5fce5ee05e095d425c8a5beb5b765b455b735c195d4b5f13616e6447677a6ad5",
      INITP_00 => X"555555aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
      INITP_01 => X"aaaaaaaaaaaaaaaaaaa955555555555555555555555555555555555555555555",
      INITP_02 => X"555555555aa5555aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
      INITP_03 => X"aaaaaaaaaaaaaaaaaaaaaaaaaa55555555555555555555555555555555555555",
      INITP_04 => X"555555aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
      INITP_05 => X"aaaaaaaaaaaaaaaaaaa955555555555555555555555555555555555555555555",
      INITP_06 => X"55555555aaaaaaaaaaaa96aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
      INITP_07 => X"aaaaaaaaaaaaaaaaaaaaaaaaaaa5555555555555555555555555555555555555",
      WRITE_MODE => "WRITE_FIRST")
   port map (
      DO   => do ( 15 downto 0),   -- 16-bit Data Output
      DOP  => do ( 17 downto 16),  -- 2-bit parity Output
      ADDR => addr (9 downto 0), -- 10-bit Address Input
      CLK  => clk,  -- Clock
      DI   => (others => '0'),   -- 8-bit Data Input
      DIP  => (others => '0'),  -- 1-bit parity Input
      EN   => '1',   -- RAM Enable Input
      SSR  => '0',  -- Synchronous Set/Reset Input
      WE   => '0'    -- Write Enable Input
   );
end behav;