library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity freqtable is
port(
	 clk : in std_logic;
	 addr : in std_logic_vector (9 downto 0);
	 en :in std_logic;
	 do : out std_logic_vector ( 17 downto 0));	 
end freqtable;

architecture Behavioral of freqtable is

begin
notes : RAMB16_S18 -- The 127 constants of how far to advance the saveform each 1/48,000th of a second
   generic map (
      INIT => X"000",
      SRVAL => X"000",
      INIT_00 => X"0064006300630062006100600060005f005e005e005d005c005c005b005a005a",
      INIT_01 => X"0070006f006f006e006d006c006b006b006a0069006800680067006600650065",
      INIT_02 => X"007e007d007c007b007a00790079007800770076007500740073007300720071",
      INIT_03 => X"008d008c008b008a00890088008700860085008400830082008200810080007f",
      INIT_04 => X"009e009d009c009b009a009900980097009600950093009200910090008f008e",
      INIT_05 => X"00b200b100af00ae00ad00ac00aa00a900a800a700a500a400a300a200a100a0",
      INIT_06 => X"00c800c600c500c300c200c000bf00be00bc00bb00ba00b800b700b600b400b3",
      INIT_07 => X"00e000de00dd00db00da00d800d600d500d300d200d000cf00cd00cc00ca00c9",
      INIT_08 => X"00fb00f900f800f600f400f200f100ef00ed00eb00ea00e800e600e500e300e2",
      INIT_09 => X"011a01180116011401120110010e010c010a0108010601040103010100ff00fd",
      INIT_0A => X"013c013a0138013601330131012f012d012b01290126012401220120011e011c",
      INIT_0B => X"01630161015e015c0159015701540152014f014d014a0148014601430141013f",
      INIT_0C => X"018f018c0189018601830180017e017b0178017601730170016e016b01680166",
      INIT_0D => X"01bf01bc01b901b601b301af01ac01a901a601a301a0019d019a019701940191",
      INIT_0E => X"01f601f201ef01eb01e801e401e101dd01da01d601d301d001cc01c901c601c3",
      INIT_0F => X"0233022f022b02270223021f021c021802140210020c02080205020101fd01fa",
      INIT_10 => X"02780274026f026b02660262025e025902550251024c024802440240023c0238",
      INIT_11 => X"02c602c102bc02b702b202ad02a802a3029e029902940290028b02860282027d",
      INIT_12 => X"031d03170311030c0306030002fb02f502f002eb02e502e002db02d502d002cb",
      INIT_13 => X"037e03780371036b0365035e03580352034c03460340033a0334032e03280322",
      INIT_14 => X"03ec03e403dd03d603cf03c803c103ba03b303ac03a6039f03980392038b0385",
      INIT_15 => X"0466045e0456044e0446043e0437042f04270420041804100409040203fa03f3",
      INIT_16 => X"04f004e704de04d504cc04c304bb04b204a904a1049804900487047f0477046f",
      INIT_17 => X"058b05810577056d05630559054f0545053b05320528051f0515050c050304f9",
      INIT_18 => X"0639062d06220617060b060005f505ea05df05d505ca05bf05b505aa05a00595",
      INIT_19 => X"06fc06ef06e206d506c906bc06b006a40697068b067f06730667065c06500644",
      INIT_1A => X"07d707c807ba07ac079e078f0782077407660758074b073d0730072307160709",
      INIT_1B => X"08cc08bc08ac089c088c087c086d085d084e083f082f08200811080307f407e5",
      INIT_1C => X"09e009ce09bc09aa0998098609750963095209410930091f090e08fe08ed08dd",
      INIT_1D => X"0b160b010aed0ad90ac50ab10a9d0a8a0a760a630a500a3d0a2a0a170a0509f2",
      INIT_1E => X"0c710c5a0c430c2d0c160c000bea0bd40bbe0ba90b930b7e0b690b540b3f0b2a",
      INIT_1F => X"0df70ddd0dc40daa0d910d780d5f0d470d2e0d160cfe0ce60cce0cb70c9f0c88",
      INIT_20 => X"0fad0f900f730f570f3b0f1e0f030ee70ecc0eb00e950e7a0e600e450e2b0e11",
      INIT_21 => X"1198117811581138111810f810d910ba109b107d105e1040102210050fe70fca",
      INIT_22 => X"13c0139b137713531330130c12e912c612a41282125f123e121c11fb11da11b9",
      INIT_23 => X"162b160215d915b115891561153a151314ec14c6149f14791454142e140913e4",
      INIT_24 => X"18e218b418861859182c180017d417a8177c1751172616fb16d116a7167d1654",
      INIT_25 => X"1bee1bba1b871b541b221af01abe1a8d1a5c1a2c19fc19cc199c196d193e1910",
      INIT_26 => X"1f591f1f1ee61ead1e751e3c1e051dce1d971d601d2a1cf41cbf1c8a1c561c21",
      INIT_27 => X"233022ef22af226f222f21f021b22174213620f920bc2080204420091fce1f93",
      INIT_28 => X"277f273626ee26a6265f261825d2258c2547250324be247b243823f523b32371",
      INIT_29 => X"2c552c032bb22b622b122ac22a742a2629d8298b293e28f228a7285c281227c8",
      INIT_2A => X"31c33167310c30b230582fff2fa72f4f2ef82ea12e4b2df62da12d4d2cfa2ca7",
      INIT_2B => X"37db3774370e36a8364435e0357c351a34b8345733f73397333832da327c321f",
      INIT_2C => X"3eb23e3e3dcb3d5a3ce93c783c093b9b3b2d3ac03a5439e8397e391438ab3842",
      INIT_2D => X"465f45dd455d44dd445e43e0436342e7426c41f2417840ff408840113f9b3f26",
      INIT_2E => X"4efd4e6c4ddb4d4c4cbd4c304ba44b184a8e4a05497c48f5486f47e9476546e1",
      INIT_2F => X"58a95806576456c35623558454e7544b53af5315527c51e4514d50b850234f90",
      INIT_30 => X"638562cd6217616360af5ffd5f4d5e9d5def5d425c965bec5b425a9a59f3594e",
      INIT_31 => X"6fb56ee76e1b6d506c876bbf6af86a33697068ad67ed672d666f65b364f7643d",
      INIT_32 => X"7d637c7c7b967ab379d178f0781277357659757f74a773d072fb722771557084",
      INIT_33 => X"8cbd8bba8ab989b988bc87c086c685ce84d783e382f081fe810f80217f357e4b",
      INIT_34 => X"9df99cd79bb69a97997a986097479630951c940992f891ea90dd8fd28ec98dc2",
      INIT_35 => X"b152b00baec7ad85ac46ab08a9cda895a75ea62aa4f8a3c8a29aa16fa0469f1f",
      INIT_36 => X"c709c59ac42ec2c5c15ebffabe99bd3abbddba83b92cb7d7b684b534b3e6b29b",
      INIT_37 => X"df69ddcddc35da9fd90dd77dd5f0d466d2dfd15acfd9ce5accdecb65c9eec87a",
      INIT_38 => X"fac5f8f7f72cf565f3a1f1e0f023ee69ecb1eafee94de79fe5f5e44de2a9e107",
      INIT_39 => X"197a17741571137211770f7f0d8b0b9b09ae07c505df03fc021e0042fe6afc96",
      INIT_3A => X"3bf239ad376b352d32f430bf2e8d2c602a37281225f023d321ba1fa41d921b84",
      INIT_3B => X"62a360165d8e5b0a588b5610539a51294ebc4c5349ef4790453442de408b3e3d",
      INIT_3C => X"8e118b34885c858a82bc7ff47d317a7377ba750672576fad6d086a6767cc6535",
      INIT_3D => X"bed1bb9ab869b53eb219aef9abdfa8cba5bda2b49fb19cb399bb96c993dc90f4",
      INIT_3E => X"f589f1edee58eac9e741e3c0e045dcd1d962d5fbd299cf3ecbe9c899c551c20e",
      INIT_3F => X"32f42ee72ae226e422ed1efe1b161735135b0f890bbd07f8043b0084fcd4f92b",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"aaaaaaa555555555555555555555555555555555555555555555555000000000",
      WRITE_MODE => "WRITE_FIRST")
   port map (
      DO   => do(15 downto 0),   -- 16-bit Data Output
      DOP  => do(17 downto 16),  -- 2-bit parity Output
      ADDR => addr, -- 10-bit Address Input
      CLK  => clk,             -- Clock
      DI   => (others => '0'),   -- 8-bit Data Input
      DIP  => (others => '0'),   -- 1-bit parity Input
      EN   => '1',               -- RAM Enable Input
      SSR  => '0',                 -- Synchronous Set/Reset Input
      WE   => '0'                -- Write Enable Input
   );
	
end Behavioral;

